library ieee;
use ieee.std_logic_1164.all;

entity MUX_3 is
	generic(g_bits:integer:=4);
	port(control:in std_logic_vector(1 downto 0);
	input0:in std_logic_vector(g_bits-1 downto 0);
	input1:in std_logic_vector(g_bits-1 downto 0);
	input2:in std_logic_vector(g_bits-1 downto 0);
	output:out std_logic_vector(g_bits-1 downto 0));
	end MUX_3;
	
Architecture MUX of MUX_3 is
begin
	process(control,input0,input1)
	begin
		case control is
			when "00"=>
				output<=input0;
			when "01"=>
				output<=input1;
			when "10"=>
				output<=input2;
			when "11"=>
				output<=(others=>'0');
			when others=>
				NULL;
			end case;
		end process;
	end MUX;